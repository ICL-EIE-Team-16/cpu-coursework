module hazard_detector(
    input logic[31:0] instruction,
    output logic hazard
);
    
endmodule